library verilog;
use verilog.vl_types.all;
entity number_analyzer_tb is
end number_analyzer_tb;
